LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.all;
USE IEEE.STD_LOGIC_UNSIGNED.all;

ENTITY keyBuffers IS
    PORT (
        clk: IN STD_LOGIC; -- master syncronos clock
        par2serLatchOut: OUT STD_LOGIC; -- 
        par2serClkOut: OUT STD_LOGIC; --
        mClear: IN STD_LOGIC; -- master clear
        shiftInA: IN STD_LOGIC; -- serial data input A
        shiftInB: IN STD_LOGIC; -- serial data input B
        
        extFifoReset: OUT STD_LOGIC; -- used to reset the external FIFO
        --extFifoFullIn: IN STD_LOGIC; -- input to tell if the FIFO is full
        extFifoWr: OUT STD_LOGIC; -- output used for write to  FIFO
        extFifoDataOut: OUT STD_LOGIC_VECTOR(14 downto 0); -- keyNumber, keyVelocity, keyState
        timerEnableOut: OUT STD_LOGIC
    );
END keyBuffers;

ARCHITECTURE keyBuffers_arch OF keyBuffers IS
    SIGNAL keyIndex: STD_LOGIC_VECTOR(6 downto 0);
    --SIGNAL keyIndex: STD_LOGIC_VECTOR(1 downto 0); -- debug
    SUBTYPE timerValue_width IS STD_LOGIC_VECTOR(6 downto 0);
    TYPE timerValue_length IS ARRAY (87 DOWNTO 0) OF timerValue_width;
    --TYPE timerValue_length IS ARRAY (3 DOWNTO 0) OF timerValue_width; -- debug
    SIGNAL timerValue: timerValue_length;

BEGIN PROCESS (clk, mClear, shiftInA, shiftInB, timerValue, keyIndex )
    variable timerEnable: STD_LOGIC;
    variable timerValueTemp: STD_LOGIC_VECTOR(6 downto 0);
    variable seqState: STD_LOGIC; --_VECTOR(1 downto 0); -- sequence state
    variable masterReset: STD_LOGIC;

    BEGIN          
        timerEnable := shiftInA and (not shiftInB);
        extFifoReset <= masterReset;
        if (clk'EVENT and clk = '1' and mClear = '1') then
            masterReset := '1';
        elsif (clk'EVENT and clk = '1' and mClear = '0') then
            masterReset := '0';
        end if;
        
        if (masterReset = '1') then
            for i in 87 downto 0 loop 
            --for i in 3 downto 0 loop -- debug
                timerValue(i) <= "0000000";
            end loop;
            keyIndex <= "1010111"; -- set to index 87 at reset
            --keyIndex <= "11"; -- debug
            seqState := '1'; -- to make par2ser latch work after an master reset
            extFifoWr <= '0'; -- active high 
            par2serLatchOut <= '1'; -- active low (on negative edge)
            par2serClkOut <= '0'; -- active high (on positive edge)
        elsif (clk'EVENT and clk = '0' and seqState = '0') then
            
            seqState := '1';
            par2serLatchOut <= '1'; -- deactivate par2ser latch (active low)
        
        elsif (clk'EVENT and clk = '0' and seqState = '1') then
            
            seqState := '0';
            if (keyIndex /= 87) then
                keyIndex <= keyIndex + "0000001";
            else
                keyIndex <= "0000000";
                par2serLatchOut <= '0'; -- (active low) fetch all keys
            end if;    
            
            timerValue(0) <= timerValueTemp;
            timerValue(87 downto 1) <= timerValue(86 downto 0);
            
        elsif (clk'EVENT and clk = '1' and seqState = '0') then 
            
            if (timerEnable = '0' and timerValue(87) /= 0) then -- write value to FIFO
                extFifoWr <= '1'; -- active high
            end if;
            par2serClkOut <= '0';
            
            if (timerEnable = '1' and timerValue(87) /= "1111111") then
                timerValueTemp := timerValue(87) + "0000001";
            elsif (timerEnable = '1') then
                timerValueTemp := "1111111";
            elsif (timerEnable = '0') then
                timerValueTemp := "0000000";
            end if;

        elsif (clk'EVENT and clk = '1' and seqState = '1') then

            par2serClkOut <= '1'; -- clock in next key'
            extFifoWr <= '0'; -- active high

        END If;
		timerEnableOut <= timerEnable;
        extFifoDataOut(14) <= shiftInA and shiftInB;
        extFifoDataOut(13 downto 7) <= keyIndex(6 downto 0);
        extFifoDataOut(6 downto 0) <= timerValue(87)(6 downto 0);
    END PROCESS;
END keyBuffers_arch;